
module FIFO(FIFO_if.DUT f1);
 
localparam max_fifo_addr = $clog2(f1.FIFO_DEPTH);

reg [f1.FIFO_WIDTH-1:0] mem [f1.FIFO_DEPTH-1:0];

reg [max_fifo_addr-1:0] wr_ptr, rd_ptr;
reg [max_fifo_addr:0] count;

always @(posedge f1.clk or negedge f1.rst_n) begin
	if (!f1.rst_n) begin
		wr_ptr <= 0;
		f1.wr_ack <= 0;
		f1.overflow <= 0;
	end
	else if (f1.wr_en && count < f1.FIFO_DEPTH) begin
		mem[wr_ptr] <= f1.data_in;
		f1.wr_ack <= 1;
		wr_ptr <= wr_ptr + 1;
	end
	else begin 
		f1.wr_ack <= 0; 
		if (f1.full & f1.wr_en)
			f1.overflow <= 1;
		else
			f1.overflow <= 0;
	end
end

always @(posedge f1.clk or negedge f1.rst_n) begin
	if (!f1.rst_n) begin
		rd_ptr <= 0;
		f1.data_out <= 0;
		f1.underflow <= 0;
	end
	else if (f1.rd_en && count != 0) begin
		f1.data_out <= mem[rd_ptr];
		rd_ptr <= rd_ptr + 1;
	end

	else begin 
		
		if (f1.empty & f1.rd_en)
			f1.underflow <= 1;
		else
			f1.underflow <= 0;
	end

end

always @(posedge f1.clk or negedge f1.rst_n) begin
	if (!f1.rst_n) begin
		count <= 0;
	end
	else begin
		if	( ({f1.wr_en, f1.rd_en} == 2'b10) && !f1.full) 
			count <= count + 1;
		else if ( ({f1.wr_en, f1.rd_en} == 2'b01) && !f1.empty)
			count <= count - 1;
			else if ( ({f1.wr_en, f1.rd_en} == 2'b11) && f1.empty)
			count <= count + 1;
			else if ( ({f1.wr_en, f1.rd_en} == 2'b11) && f1.full)
			count <= count - 1;
			
	end
end

assign f1.full = (count == f1.FIFO_DEPTH)? 1 : 0;
assign f1.empty = (count == 0)? 1 : 0;
assign f1.almostfull = (count == f1.FIFO_DEPTH-1)? 1 : 0; 
assign f1.almostempty = (count == 1)? 1 : 0;

`ifdef SIM


always_comb begin 
    if (!f1.rst_n) begin
       p1:assert final(f1.full == 0 && f1.empty == 1 && f1.almostfull == 0 && f1.almostempty == 0 && 
	   f1.underflow == 0 && f1.overflow == 0 && f1.wr_ack == 0 && rd_ptr == 0 && wr_ptr == 0 && count == 0);
    end
end


property p2;
@(posedge f1.clk) disable iff (!f1.rst_n) (f1.wr_en && !f1.full) |-> ##1 (f1.wr_ack == 1);
endproperty

assert property (p2); 
cover property (p2);


property p3;
@(posedge f1.clk) disable iff (!f1.rst_n) (f1.wr_en && f1.full) |-> ##1 (f1.overflow == 1);
endproperty

assert property (p3); 
cover property (p3);


property p4;
@(posedge f1.clk) disable iff (!f1.rst_n) (f1.rd_en && f1.empty) |-> ##1 (f1.underflow == 1);
endproperty

assert property (p4); 
cover property (p4);


property p5;
@(posedge f1.clk) disable iff (!f1.rst_n) (count == 0) |-> (f1.empty == 1);
endproperty

assert property (p5); 
cover property (p5);


property p6;
@(posedge f1.clk) disable iff (!f1.rst_n) (count == f1.FIFO_DEPTH) |-> (f1.full == 1);
endproperty

assert property (p6); 
cover property (p6);


property p7;
@(posedge f1.clk) disable iff (!f1.rst_n) (count == (f1.FIFO_DEPTH - 'b1)) |-> (f1.almostfull == 1);
endproperty

assert property (p7); 
cover property (p7);

property p8;
@(posedge f1.clk) disable iff (!f1.rst_n) (count == 1) |-> (f1.almostempty == 1);
endproperty

assert property (p8); 
cover property (p8);


property p9;
@(posedge f1.clk) disable iff (!f1.rst_n) ((!f1.rd_en throughout f1.wr_en[->8]) ##0 (wr_ptr == 0)) |-> (wr_ptr == 0);
endproperty

assert property (p9); 
cover property (p9);


property p10;
@(posedge f1.clk) disable iff (!f1.rst_n) ((!f1.wr_en throughout f1.rd_en[->8]) ##0 (rd_ptr == 0)) |-> (rd_ptr == 0);
endproperty

assert property (p10); 
cover property (p10);

always @(posedge f1.clk) begin
	p11:assert final(rd_ptr < (f1.FIFO_DEPTH) && wr_ptr < (f1.FIFO_DEPTH) && count <= (f1.FIFO_DEPTH));
end

`endif 
endmodule




